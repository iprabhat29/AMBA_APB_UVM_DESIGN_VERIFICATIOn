package mypackage;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "my_config.svh"
	`include "mytransaction.svh"
	`include "mysequencer.svh"
	`include "mydriver.svh"
	`include "myagent.svh"	
endpackage